module part1 (SW, LEDR, HEX1, HEX0);
	input [7:0] SW;
	output [7:0] LEDR;
	output [6:0] HEX1, HEX0;

	//LED to switch
	assign LEDR = SW;
	
	//SW[7:4]
	assign HEX1 = (SW[7:4] == 4'b1001) ? 7'b0010000 : 
                  (SW[7:4] == 4'b1000) ? 7'b0000000 : 
                  (SW[7:4] == 4'b0111) ? 7'b1111000 : 
                  (SW[7:4] == 4'b0110) ? 7'b0000010 : 
                  (SW[7:4] == 4'b0101) ? 7'b0010010 : 
                  (SW[7:4] == 4'b0100) ? 7'b0011001 : 
                  (SW[7:4] == 4'b0011) ? 7'b0110000 : 
                  (SW[7:4] == 4'b0010) ? 7'b0100100 : 
                  (SW[7:4] == 4'b0001) ? 7'b1111001 : 
                  (SW[7:4] == 4'b0000) ? 7'b1000000 : 
                  7'b1111111; // Empty
	
	//SW[7:4]
	assign HEX0 = (SW[3:0] == 4'b1001) ? 7'b0010000 : 
                  (SW[3:0] == 4'b1000) ? 7'b0000000 : 
                  (SW[3:0] == 4'b0111) ? 7'b1111000 : 
                  (SW[3:0] == 4'b0110) ? 7'b0000010 : 
                  (SW[3:0] == 4'b0101) ? 7'b0010010 : 
                  (SW[3:0] == 4'b0100) ? 7'b0011001 : 
                  (SW[3:0] == 4'b0011) ? 7'b0110000 : 
                  (SW[3:0] == 4'b0010) ? 7'b0100100 : 
                  (SW[3:0] == 4'b0001) ? 7'b1111001 : 
                  (SW[3:0] == 4'b0000) ? 7'b1000000 : 
                  7'b1111111; // Empty
	
endmodule
