module part2 (SW, HEX1, HEX0);
    input [3:0] SW;
    output [6:0] HEX1, HEX0;

    wire z;
    wire [3:0] A;

    assign z = (SW > 4'b1001);

    assign A = (SW == 4'b1010) ? 4'b0000 :
               (SW == 4'b1011) ? 4'b0001 :
               (SW == 4'b1100) ? 4'b0010 :
               (SW == 4'b1101) ? 4'b0011 :
               (SW == 4'b1110) ? 4'b0100 :
               (SW == 4'b1111) ? 4'b0101 :
               4'b0000; // Default

    wire [3:0] d0 = z ? A : SW;

    assign HEX1 = z ? 7'b1111001 : 7'b1000000;

    assign HEX0 = (d0 == 4'b1001) ? 7'b0010000 : 
                  (d0 == 4'b1000) ? 7'b0000000 :
                  (d0 == 4'b0111) ? 7'b1111000 :
                  (d0 == 4'b0110) ? 7'b0000010 :
                  (d0 == 4'b0101) ? 7'b0010010 : 
                  (d0 == 4'b0100) ? 7'b0011001 :
                  (d0 == 4'b0011) ? 7'b0110000 :
                  (d0 == 4'b0010) ? 7'b0100100 :
                  (d0 == 4'b0001) ? 7'b1111001 :
                  (d0 == 4'b0000) ? 7'b1000000 :
                  7'b1111111;
endmodule